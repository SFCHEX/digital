module add_sub_signal(input reverse,signal, output add, sub);
    wire reverse_i;
    not(reverese_i,revere)
    and(add,reverse_i,signal);
    and(sub,reverse,signal)
endmodule