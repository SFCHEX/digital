module m3216(input [15:0]i0,i1,input s,output [15:0]out)

m21 m0(out[0],i0[0],i1[0],s)
m21 m1(out[1],i0[1],i1[1],s)
m21 m2(out[2],i0[2],i1[2],s)
m21 m3(out[3],i0[3],i1[3],s)
m21 m0(out[4],i0[4],i1[4],s)
m21 m0(out[5],i0[5],i1[5],s)
m21 m0(out[6],i0[6],i1[6],s)
m21 m0(out[7],i0[7],i1[7],s)
m21 m0(out[8],i0[8],i1[8],s)
m21 m0(out[9],i0[9],i1[9],s)
m21 m0(out[10],i0[10],i1[10],s)
m21 m0(out[11],i0[11],i1[11],s)
m21 m0(out[12],i0[12],i1[12],s)
m21 m0(out[13],i0[13],i1[13],s)
m21 m0(out[14],i0[14],i1[14],s)
m21 m0(out[15],i0[15],i1[15],s)

endmodule